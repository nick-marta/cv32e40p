//////////////////////
// TODO remove
//////////////////////
module hvl_top;
  import uvm_pkg::*;
  import alu_pkg::*;
  
  initial run_test();
endmodule
